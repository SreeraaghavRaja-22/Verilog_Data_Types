module adder_tree(
    input [3:0] a, 
    input [3:]
)