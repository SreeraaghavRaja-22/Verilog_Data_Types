module encoder 8to3(
    input [7:0] d, 
    
)