module conditional_operator(); 

    integer result; 
    integer a = 9; 
    integer b = 32; 
    integer c = 0; 

    initial begin 
        #1; result = (a == 9) ? 1 : 0; 
        $display("result = %0d", result);

        #1; result = ((a + b) == 40) ? 1 : 0; 
        $display("result = %0d", result);

        #1; result = (b == 30) ? 679 : -99; 
        $display("result = %0d", result);

        #1; result = (b == 32) ? 1'bZ : 1'b0;
        $display("result = %0d", result);
        #1; 
    end 

endmodule